module alternate_debouncing_circuit  

(
    
);

endmodule //alternate_debouncing_circuit